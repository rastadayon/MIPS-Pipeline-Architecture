module cu(input [5:0] opcode, function, output Rtype, lw, sw, j , beq, bne, pcSrc, memWrite, memRead, ALUsrc, regDest, regWrite, memToReg,  output [2:0] ALUop);
endmodule
